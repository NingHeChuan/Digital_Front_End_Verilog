module foo(/*AUTOARG*/
   // Outputs
   o,
   // Inputs
   i
   );

input i;
output [DWIDTH-1:0] o;

endmodule
